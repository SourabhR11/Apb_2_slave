                                	             		     		     		     	             		     		     		     		     	             		     		     	             	             	             		     		     	                                 endmodule
