`include "uvm_macros.svh"
import uvm_pkg::*;

//`include "apb_design.sv"
`include "defines.svh"
`include "apb_intf.sv"
`include "apb_seq_item.sv"
`include "apb_seq.sv"
`include "apb_seqr.sv"
`include "apb_driver.sv"
`include "apb_ip_mon.sv"
`include "apb_op_mon.sv"
`include "apb_active_agent.sv"
`include "apb_passive_agent.sv"
`include "apb_sb.sv"
`include "apb_cov.sv"
`include "apb_env.sv"
`include "apb_test.sv"
